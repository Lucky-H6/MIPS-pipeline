module Instruction_Memory(ReadAddr, Ins);

    input [31:0] ReadAddr;
    output reg [31:0] Ins;

    always @(*) begin
        if (ReadAddr == 32'h80000004)
            Ins <= 32'h0810008e;
        else
            case ({1'b0, ReadAddr[30:0]})
                32'h00400004: Ins <= 32'h3c014000;
                32'h00400008: Ins <= 32'h34280000;
                32'h0040000C: Ins <= 32'had000008;
                32'h00400010: Ins <= 32'h240b6d60;
                32'h00400014: Ins <= 32'h240a0000;
                32'h00400018: Ins <= 32'had0b0000;
                32'h0040001C: Ins <= 32'had0a0004;
                32'h00400020: Ins <= 32'h240b0003;
                32'h00400024: Ins <= 32'had0b0008;
                32'h00400028: Ins <= 32'h3c014000;
                32'h0040002C: Ins <= 32'h34290014;
                32'h00400030: Ins <= 32'h8d3b0000;
                32'h00400034: Ins <= 32'h24100000;
                32'h00400038: Ins <= 32'h2411007f;
                32'h0040003C: Ins <= 32'h00102021;
                32'h00400040: Ins <= 32'h24050000;
                32'h00400044: Ins <= 32'h00113021;
                32'h00400048: Ins <= 32'h0c100015;
                32'h0040004C: Ins <= 32'h00000000;
                32'h00400050: Ins <= 32'h081000f4;
                32'h00400054: Ins <= 32'h23bdffe4;
                32'h00400058: Ins <= 32'hafb50018;
                32'h0040005C: Ins <= 32'hafb40014;
                32'h00400060: Ins <= 32'hafb30010;
                32'h00400064: Ins <= 32'hafb2000c;
                32'h00400068: Ins <= 32'hafb10008;
                32'h0040006C: Ins <= 32'hafb00004;
                32'h00400070: Ins <= 32'hafbf0000;
                32'h00400074: Ins <= 32'h00048021;
                32'h00400078: Ins <= 32'h00058821;
                32'h0040007C: Ins <= 32'h00069021;
                32'h00400080: Ins <= 32'h0005a021;
                32'h00400084: Ins <= 32'h0006a821;
                32'h00400088: Ins <= 32'h00144080;
                32'h0040008C: Ins <= 32'h01104020;
                32'h00400090: Ins <= 32'h8d130000;
                32'h00400094: Ins <= 32'h00124080;
                32'h00400098: Ins <= 32'h01104020;
                32'h0040009C: Ins <= 32'h8d080000;
                32'h004000A0: Ins <= 32'h00000000;
                32'h004000A4: Ins <= 32'h0113402a;
                32'h004000A8: Ins <= 32'h34010001;
                32'h004000AC: Ins <= 32'h00284023;
                32'h004000B0: Ins <= 32'h0232482a;
                32'h004000B4: Ins <= 32'h01094024;
                32'h004000B8: Ins <= 32'h00000000;
                32'h004000BC: Ins <= 32'h1100000c;
                32'h004000C0: Ins <= 32'h2252ffff;
                32'h004000C4: Ins <= 32'h00124080;
                32'h004000C8: Ins <= 32'h01104020;
                32'h004000CC: Ins <= 32'h8d080000;
                32'h004000D0: Ins <= 32'h00000000;
                32'h004000D4: Ins <= 32'h0113402a;
                32'h004000D8: Ins <= 32'h34010001;
                32'h004000DC: Ins <= 32'h00284023;
                32'h004000E0: Ins <= 32'h0232482a;
                32'h004000E4: Ins <= 32'h01094024;
                32'h004000E8: Ins <= 32'h00000000;
                32'h004000EC: Ins <= 32'h1500fff4;
                32'h004000F0: Ins <= 32'h00114080;
                32'h004000F4: Ins <= 32'h01104020;
                32'h004000F8: Ins <= 32'h8d080000;
                32'h004000FC: Ins <= 32'h00000000;
                32'h00400100: Ins <= 32'h0268402a;
                32'h00400104: Ins <= 32'h34010001;
                32'h00400108: Ins <= 32'h00284023;
                32'h0040010C: Ins <= 32'h0232482a;
                32'h00400110: Ins <= 32'h01094024;
                32'h00400114: Ins <= 32'h00000000;
                32'h00400118: Ins <= 32'h1100000c;
                32'h0040011C: Ins <= 32'h22310001;
                32'h00400120: Ins <= 32'h00114080;
                32'h00400124: Ins <= 32'h01104020;
                32'h00400128: Ins <= 32'h8d080000;
                32'h0040012C: Ins <= 32'h00000000;
                32'h00400130: Ins <= 32'h0268402a;
                32'h00400134: Ins <= 32'h34010001;
                32'h00400138: Ins <= 32'h00284023;
                32'h0040013C: Ins <= 32'h0232482a;
                32'h00400140: Ins <= 32'h01094024;
                32'h00400144: Ins <= 32'h00000000;
                32'h00400148: Ins <= 32'h1500fff4;
                32'h0040014C: Ins <= 32'h0232402a;
                32'h00400150: Ins <= 32'h00000000;
                32'h00400154: Ins <= 32'h15000002;
                32'h00400158: Ins <= 32'h08100060;
                32'h0040015C: Ins <= 32'h00000000;
                32'h00400160: Ins <= 32'h00112080;
                32'h00400164: Ins <= 32'h00122880;
                32'h00400168: Ins <= 32'h02042020;
                32'h0040016C: Ins <= 32'h02052820;
                32'h00400170: Ins <= 32'h0c100088;
                32'h00400174: Ins <= 32'h00000000;
                32'h00400178: Ins <= 32'h08100025;
                32'h0040017C: Ins <= 32'h00000000;
                32'h00400180: Ins <= 32'h00144080;
                32'h00400184: Ins <= 32'h02084020;
                32'h00400188: Ins <= 32'h00114880;
                32'h0040018C: Ins <= 32'h02094820;
                32'h00400190: Ins <= 32'h8d290000;
                32'h00400194: Ins <= 32'h00000000;
                32'h00400198: Ins <= 32'had090000;
                32'h0040019C: Ins <= 32'h00114080;
                32'h004001A0: Ins <= 32'h02084020;
                32'h004001A4: Ins <= 32'had130000;
                32'h004001A8: Ins <= 32'h2228ffff;
                32'h004001AC: Ins <= 32'h0288402a;
                32'h004001B0: Ins <= 32'h00000000;
                32'h004001B4: Ins <= 32'h11000005;
                32'h004001B8: Ins <= 32'h00102021;
                32'h004001BC: Ins <= 32'h00142821;
                32'h004001C0: Ins <= 32'h2226ffff;
                32'h004001C4: Ins <= 32'h0c100015;
                32'h004001C8: Ins <= 32'h00000000;
                32'h004001CC: Ins <= 32'h22280001;
                32'h004001D0: Ins <= 32'h0115402a;
                32'h004001D4: Ins <= 32'h00000000;
                32'h004001D8: Ins <= 32'h11000005;
                32'h004001DC: Ins <= 32'h00102021;
                32'h004001E0: Ins <= 32'h22250001;
                32'h004001E4: Ins <= 32'h00153021;
                32'h004001E8: Ins <= 32'h0c100015;
                32'h004001EC: Ins <= 32'h00000000;
                32'h004001F0: Ins <= 32'h00001020;
                32'h004001F4: Ins <= 32'h8fb50018;
                32'h004001F8: Ins <= 32'h8fb40014;
                32'h004001FC: Ins <= 32'h8fb30010;
                32'h00400200: Ins <= 32'h8fb2000c;
                32'h00400204: Ins <= 32'h8fb10008;
                32'h00400208: Ins <= 32'h8fb00004;
                32'h0040020C: Ins <= 32'h8fbf0000;
                32'h00400210: Ins <= 32'h23bd001c;
                32'h00400214: Ins <= 32'h00000000;
                32'h00400218: Ins <= 32'h03e00008;
                32'h0040021C: Ins <= 32'h00000000;
                32'h00400220: Ins <= 32'h8c880000;
                32'h00400224: Ins <= 32'h8ca90000;
                32'h00400228: Ins <= 32'haca80000;
                32'h0040022C: Ins <= 32'hac890000;
                32'h00400230: Ins <= 32'h03e00008;
                32'h00400234: Ins <= 32'h00000000;
                32'h00400238: Ins <= 32'h2408000f;
                32'h0040023C: Ins <= 32'h013bd824;
                32'h00400240: Ins <= 32'h24080000;
                32'h00400244: Ins <= 32'h00000000;
                32'h00400248: Ins <= 32'h1368002d;
                32'h0040024C: Ins <= 32'h24080001;
                32'h00400250: Ins <= 32'h00000000;
                32'h00400254: Ins <= 32'h1368002d;
                32'h00400258: Ins <= 32'h24080002;
                32'h0040025C: Ins <= 32'h00000000;
                32'h00400260: Ins <= 32'h1368002d;
                32'h00400264: Ins <= 32'h24080003;
                32'h00400268: Ins <= 32'h00000000;
                32'h0040026C: Ins <= 32'h1368002d;
                32'h00400270: Ins <= 32'h24080004;
                32'h00400274: Ins <= 32'h00000000;
                32'h00400278: Ins <= 32'h1368002d;
                32'h0040027C: Ins <= 32'h24080005;
                32'h00400280: Ins <= 32'h00000000;
                32'h00400284: Ins <= 32'h1368002d;
                32'h00400288: Ins <= 32'h24080006;
                32'h0040028C: Ins <= 32'h00000000;
                32'h00400290: Ins <= 32'h1368002d;
                32'h00400294: Ins <= 32'h24080007;
                32'h00400298: Ins <= 32'h00000000;
                32'h0040029C: Ins <= 32'h1368002d;
                32'h004002A0: Ins <= 32'h24080008;
                32'h004002A4: Ins <= 32'h00000000;
                32'h004002A8: Ins <= 32'h1368002d;
                32'h004002AC: Ins <= 32'h24080009;
                32'h004002B0: Ins <= 32'h00000000;
                32'h004002B4: Ins <= 32'h1368002d;
                32'h004002B8: Ins <= 32'h2408000a;
                32'h004002BC: Ins <= 32'h00000000;
                32'h004002C0: Ins <= 32'h1368002d;
                32'h004002C4: Ins <= 32'h2408000b;
                32'h004002C8: Ins <= 32'h00000000;
                32'h004002CC: Ins <= 32'h1368002d;
                32'h004002D0: Ins <= 32'h2408000c;
                32'h004002D4: Ins <= 32'h00000000;
                32'h004002D8: Ins <= 32'h1368002d;
                32'h004002DC: Ins <= 32'h2408000d;
                32'h004002E0: Ins <= 32'h00000000;
                32'h004002E4: Ins <= 32'h1368002d;
                32'h004002E8: Ins <= 32'h2408000e;
                32'h004002EC: Ins <= 32'h00000000;
                32'h004002F0: Ins <= 32'h1368002d;
                32'h004002F4: Ins <= 32'h2408000f;
                32'h004002F8: Ins <= 32'h00000000;
                32'h004002FC: Ins <= 32'h1368002d;
                32'h00400300: Ins <= 32'h240901fc;
                32'h00400304: Ins <= 32'h081000f0;
                32'h00400308: Ins <= 32'h00000000;
                32'h0040030C: Ins <= 32'h24090160;
                32'h00400310: Ins <= 32'h081000f0;
                32'h00400314: Ins <= 32'h00000000;
                32'h00400318: Ins <= 32'h240901da;
                32'h0040031C: Ins <= 32'h081000f0;
                32'h00400320: Ins <= 32'h00000000;
                32'h00400324: Ins <= 32'h240901f2;
                32'h00400328: Ins <= 32'h081000f0;
                32'h0040032C: Ins <= 32'h00000000;
                32'h00400330: Ins <= 32'h24090166;
                32'h00400334: Ins <= 32'h081000f0;
                32'h00400338: Ins <= 32'h00000000;
                32'h0040033C: Ins <= 32'h240901b6;
                32'h00400340: Ins <= 32'h081000f0;
                32'h00400344: Ins <= 32'h00000000;
                32'h00400348: Ins <= 32'h240901be;
                32'h0040034C: Ins <= 32'h081000f0;
                32'h00400350: Ins <= 32'h00000000;
                32'h00400354: Ins <= 32'h240901e0;
                32'h00400358: Ins <= 32'h081000f0;
                32'h0040035C: Ins <= 32'h00000000;
                32'h00400360: Ins <= 32'h240901fe;
                32'h00400364: Ins <= 32'h081000f0;
                32'h00400368: Ins <= 32'h00000000;
                32'h0040036C: Ins <= 32'h240901f6;
                32'h00400370: Ins <= 32'h081000f0;
                32'h00400374: Ins <= 32'h00000000;
                32'h00400378: Ins <= 32'h240901ef;
                32'h0040037C: Ins <= 32'h081000f0;
                32'h00400380: Ins <= 32'h00000000;
                32'h00400384: Ins <= 32'h240901ff;
                32'h00400388: Ins <= 32'h081000f0;
                32'h0040038C: Ins <= 32'h00000000;
                32'h00400390: Ins <= 32'h2409019d;
                32'h00400394: Ins <= 32'h081000f0;
                32'h00400398: Ins <= 32'h00000000;
                32'h0040039C: Ins <= 32'h240901fd;
                32'h004003A0: Ins <= 32'h081000f0;
                32'h004003A4: Ins <= 32'h00000000;
                32'h004003A8: Ins <= 32'h2409019f;
                32'h004003AC: Ins <= 32'h081000f0;
                32'h004003B0: Ins <= 32'h00000000;
                32'h004003B4: Ins <= 32'h2409018f;
                32'h004003B8: Ins <= 32'h081000f0;
                32'h004003BC: Ins <= 32'h00000000;
                32'h004003C0: Ins <= 32'h3c014000;
                32'h004003C4: Ins <= 32'h342a0010;
                32'h004003C8: Ins <= 32'had490000;
                32'h004003CC: Ins <= 32'h03400008;
                32'h004003D0: Ins <= 32'h3c014000;
                32'h004003D4: Ins <= 32'h34280014;
                32'h004003D8: Ins <= 32'h8d090000;
                32'h004003DC: Ins <= 32'h00000000;
                32'h004003E0: Ins <= 32'h013bd822;
                32'h80000004: Ins <= 32'h0810008e;
                default: Ins <= 32'h00000000;
        endcase
    end

endmodule